module hola (
    input wire a, // Signal de entrada de tipo wire (Se utilia para vables)
    output wire y // Es una salida de tipo wire, es un cable que transporta la señal de salida
);

endmodule
